`timescale 1ns / 1ps

module tb_convolution_top_alt;

// --- Parameters ---
parameter PIXEL_W  = 16;
parameter KERNEL_W = 16;
parameter RESULT_W = 48;
parameter IMG_SIZE = 8'd128;
parameter CHANNELS = 9'd64;

// --- Clock & Reset ---
reg clk;
reg aresetn;

// --- UUT Signals ---
reg Load_kernel_BRAM;
wire [255:0] kernel_BRAM_doutb;
wire enb_kernel_BRAM;
wire [7:0] kernel_BRAM_counter_out;
reg [47:0] bias_val;

// Slave AXI-Stream (Input)
reg [PIXEL_W-1:0] s_axis_tdata;
reg s_axis_tvalid;
wire s_axis_tready;
reg s_axis_tlast;

// Master AXI-Stream (Output)
wire [63:0] m_axis_tdata;
wire m_axis_tvalid;
reg m_axis_tready;
wire m_axis_tlast;

// --- Reference Model Memories ---
reg signed [PIXEL_W-1:0]  ref_input  [0:CHANNELS-1][0:IMG_SIZE-1][0:IMG_SIZE-1];
reg signed [KERNEL_W-1:0] ref_kernel [0:CHANNELS-1][0:2][0:2]; // 3x3 kernels
reg signed [RESULT_W-1:0] ref_output [0:IMG_SIZE-1][0:IMG_SIZE-1];

// --- Simulation Internal Variables ---
integer i, j, k, r, c, ch;
integer image_index;
integer err_count = 0;
integer pixels_received = 0;

// --- UUT Instantiation ---
convolution_top uut (
    .clk(clk),
    .aresetn(aresetn),
    .Load_kernel_BRAM(Load_kernel_BRAM),
    .Image_size(IMG_SIZE),
    .Channel_size(CHANNELS),
    .kernel_BRAM_doutb(kernel_BRAM_doutb),
    .enb_kernel_BRAM(enb_kernel_BRAM),
    .kernel_BRAM_counter_out(kernel_BRAM_counter_out),
    .bias_BRAM_douta(bias_val),
    .s_axis_tdata(s_axis_tdata),
    .s_axis_tvalid(s_axis_tvalid),
    .s_axis_tready(s_axis_tready),
    .s_axis_tlast(s_axis_tlast),
    .m_axis_tdata(m_axis_tdata),
    .m_axis_tvalid(m_axis_tvalid),
    .m_axis_tready(m_axis_tready),
    .m_axis_tlast(m_axis_tlast)
);

// --- Clock Generation ---
initial clk = 0;
always #5 clk = ~clk;

// Mock S_AXIS for image (storing one full image, all channels)
reg signed [PIXEL_W-1:0] image_mem [0:1048575];

// Kernel BRAM (storing 1 kernel)
reg signed [143:0] kernel_mem [0:CHANNELS-1];

assign kernel_BRAM_doutb = {112'b0, kernel_mem[kernel_BRAM_counter_out]};

always @(posedge clk) begin
    s_axis_tdata <= image_mem[image_index];
end

// Simulasi stimulus sinyal input
initial begin
    // Load the files generated by Python
    $readmemh("image_data_hex.mem",  image_mem);
    $readmemh("kernel_data.mem", kernel_mem);

    // Init data
    aresetn = 0;
    Load_kernel_BRAM = 0;
    s_axis_tvalid = 0;
    m_axis_tready = 1;
    bias_val = 48'd652;
    s_axis_tlast = 0;

    @(posedge clk);
    aresetn = 1;
    Load_kernel_BRAM = 0;
    s_axis_tvalid = 0;
    m_axis_tready = 1;

    @(posedge clk);
    Load_kernel_BRAM = 1;
    s_axis_tvalid = 0;
    m_axis_tready = 1;

    @(posedge clk);
    @(posedge clk);
    @(posedge clk);
    @(posedge clk);
    @(posedge clk);

    Load_kernel_BRAM = 0;
    s_axis_tvalid = 0;
    m_axis_tready = 1;

    @(posedge clk);
    s_axis_tvalid = 1;
    m_axis_tready = 1;

    @(posedge clk);
    @(posedge clk);
    @(posedge clk);
    @(posedge clk);
end

endmodule